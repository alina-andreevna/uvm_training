package tb_pkg;
    import uvm_pkg::*;

    virtual interface fir_if global_fir_if;

    `include "uvm_macros.svh"
    `include "data_seq_item.svh"
    `include "data_sequencer.svh"
    `include "data_sequence.svh"
    `include "data_driver.svh"
    `include "data_monitor.svh"
    `include "data_scoreboard.svh"
    `include "data_agent.svh"
    `include "data_env.svh"  
    `include "verbose_test.svh"
endpackage: tb_pkg
