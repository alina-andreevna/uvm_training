package fir_param_pkg;

  `define CLK_PERIOD 10ns

  `define INPUT_WORD_SIZE 10
  `define OUTPUT_WORD_SIZE 10

endpackage: fir_param_pkg