`include  "sq_base.sv"
`include  "tst_base.sv"
`include  "sq_start.sv"
`include  "tst_start.sv"