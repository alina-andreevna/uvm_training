package tb_pkg;
  import uvm_pkg::*;

  virtual interface fir_if global_fir_if;

  `include "uvm_macros.svh"
  `include "driver.svh"
  `include "scoreboard.svh"
  `include "printer.svh"
  `include "tester_env.svh"  
  `include "verbose_test.svh"
endpackage: tb_pkg
